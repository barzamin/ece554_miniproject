module tpumac_tb();
  logic clk, rst_n;
  logic en, WrEn;

  logic signed [7:0] A;
  logic signed [7:0] B;
  logic signed [15:0] C;
endmodule
